`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: SRI KRISHNA G
// 
// Create Date:    15:35:39 03/25/2023 
// Design Name: LOGICAL OR GATE
// Module Name:    OR_gate 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module OR_gate(in1,in2,out);
input in1,in2;
output out;
assign out = in1|in2;
endmodule
